* C:\Users\Tarush\eSim-Workspace\D_FF_New\D_FF_New.cir

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

xM13  CLK_BAR CLK vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM14  CLK_BAR CLK GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM1  Net-_M1-Pad1_ D_IN vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM2  Net-_C1-Pad1_ CLK Net-_M1-Pad1_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM6  Net-_C1-Pad1_ CLK_BAR Net-_M6-Pad3_ GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM7  Net-_M6-Pad3_ D_IN GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
C1  Net-_C1-Pad1_ GND 0.0001u		
xM3  Qm Net-_C1-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM8  Qm Net-_C1-Pad1_ GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM4  Net-_M4-Pad1_ Qm vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM5  Net-_C2-Pad1_ CLK_BAR Net-_M4-Pad1_ vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM9  Net-_C2-Pad1_ CLK Net-_M10-Pad1_ GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
xM10  Net-_M10-Pad1_ Qm GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		
C2  Net-_C2-Pad1_ GND 0.0001u		
xM11  Qs Net-_C2-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5		
xM12  Qs Net-_C2-Pad1_ GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5		

Vdd vdd 0 5

* pulse command(Vintial Von Tdelay Trise Tfall Ton Ttotal Ncycles)
Vd0 D_IN 0 pulse(0 5 7m 10p 10p 10m 20m)
Vd1 CLK 0 pulse(0 5 0s 10p 10p 6m 12m)

.tran 0.002ms 100ms

.control
run

plot V(CLK) V(D_IN) V(Qm) V(Qs) 

.endc		

.end
